library IEEE;
use ieee.std_logic_1164.all;

entity top_level is
  port (
    HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7 : OUT STD_LOGIC_VECTOR(6 downto 0)
  );
end entity;